module hello ();
    initial begin
        $display("\n\t Hello  World\n");
    end    
endmodule